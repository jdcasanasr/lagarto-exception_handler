package riscv_pkg;

    localparam XLEN = 64;

endpackage